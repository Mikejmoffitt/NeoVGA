-- neovga.vhd
-- NeoVGA Rev 2
-- 2015 Michael Moffitt
-------------------------
--
-- Top level entity for NeoVGA.
--
-- Neo-Geo Wiring Notes:
-- RGB pixel bus is 5 bits per channel with 0 as the LSB. Locations will
-- differ between different models.
--
-- DAK and SHAD should be pulled before the 74LS05, or else the mixed-in
-- analogue RGB levels will screw with the FPGA's ability to correctly
-- read the digital data. It is worth noting that they will be inverted.
-- That is what NeoVGA expects. The 74LS05's are open collectors so the
-- DAK and SHAD signals only pull it down when asserted.
--
-- The Neo clock is pulled from the 68000 CPU, generated by a division of
-- the master 24MHz clock. If you would like to divide this yourself then
-- by all means go ahead. I won't recommend pulling off of the 24Mhz clock
-- directly only because it often causes my Neo-Geo to reset. I have not 
-- explored this issue much so it may be a non-issue. 
--
-- The sync signal is the Neo-Geo's composite sync signal, which should be
-- pulled before it is put through a voltage divider on the JAMMA edge. 
-- The neo_clr_n signal is the blanking signal on the original DAC's '273s
-- clear input. On early MVS systems, this blanks the screen during the
-- top and bottom borders and during retrace so palette writes are not
-- seen on screen. On later systems (like MV-1C) the blanking signal is 
-- active during the horizontal front and back porch as well. 
--
-- Not all boards have the same sync timings, so adjustments may be needed
-- for different models.

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity neovga is 
generic (vga_depth: integer := 10);
port (
	-- Neo-Geo pixel bus data and timing sources
	neo_clk: in std_logic; -- Port D 0;
	neo_dak: in std_logic; -- Port D 1;
	neo_shad: in std_logic; -- Port D 2;
	neo_clr_n: in std_logic; -- Port D 3;
	neo_csync: in std_logic; -- Port D 7;
	
	-- User switches
	sw_ypbpr_n: in std_logic; -- SW1
	sw_scanlines_n: in std_logic_vector(1 downto 0); -- SW2, SW3
	sw_sdtv_res_n: in std_logic; -- SW4
	
	j_mv1c_sel_n: in std_logic; -- J1
	j_want_sog_n: in std_logic; -- J2
	
	neo_red: in std_logic_vector(4 downto 0); -- Port A 0 - 4;
	neo_green: in std_logic_vector(4 downto 0); -- Port B 0 - 4
	neo_blue: in std_logic_vector(4 downto 0); -- Port C 0 - 4
	
	led_out: out std_logic;
	
	-- VGA outputs
	vga_red: out std_logic_vector(vga_depth - 1 downto 0);
	vga_green: out std_logic_vector(vga_depth - 1 downto 0);
	vga_blue: out std_logic_vector(vga_depth - 1 downto 0);
	vga_clk: out std_logic;
	vga_blank: out std_logic;
	vga_hsync: out std_logic;
	vga_vsync: out std_logic;
	vga_sync: out std_logic
	);
end neovga;

architecture behavioral of neovga is 
constant FAKESYNC_THRESH: integer := 64;

--------- Timings for different chipset generations -----------
constant NEO_GRZ_SHIFT: integer := 24;
constant PRO_B0_SHIFT: integer := 704;
constant NEO_B1_SHIFT: integer := PRO_B0_SHIFT;
---------------------------------------------------

-- The H shift must be adjusted to match the appropriate Neo-Geo graphics
-- chipset.

-- Defaults to B0/B1 shift amount; if a GRZ (MV-1C, single-game board) is detected this will get overwritten.
signal h_shift: integer := PRO_B0_SHIFT;

-- Indeces for colors inside one 17-bit pixel packet
constant RED_POS: integer := 16;
constant GREEN_POS: integer := 11;
constant BLUE_POS: integer := 6;
constant DEPTH_BITS: integer := 5;
constant RED_END: integer := RED_POS - DEPTH_BITS + 1;
constant GREEN_END: integer := GREEN_POS - DEPTH_BITS + 1;
constant BLUE_END: integer := BLUE_POS - DEPTH_BITS + 1;

-- VGA output timings
constant VGA_VISIBLE_START: integer := 0;
constant VGA_VISIBLE_END: integer := 332;
constant VGA_HSYNC_START: integer := 332;
constant VGA_HSYNC_END: integer := 378;
constant NUM_LINES: integer := 264;
constant VGA_VSYNC_LINE_START: integer := 260;
constant VGA_VSYNC_LINE_END: integer := 262;

-- Common constants
constant U17_ZERO: std_logic_vector(16 downto 0) := "00000000000000000";
constant U16_ZERO: std_logic_vector(15 downto 0) := "0000000000000000";

-- Line length in clocks (2x Neo-Geo pixel clock, 1/2 standard 640x480 pixel clock).
constant VGA_LINE_LEN: integer := 384;
constant NEO_LINE_LEN: integer := 768;

signal vsync_count: std_logic_vector(15 downto 0) := U16_ZERO;
signal neo_pxcount: std_logic_vector(15 downto 0) := U16_ZERO;
signal vga_pxcount: std_logic_vector(15 downto 0) := U16_ZERO;
signal line_count: std_logic_vector(15 downto 0) := U16_ZERO;

-- C-sync decoding
-- Increase to shift to the right
signal fakesync_delayed: std_logic;
signal sync_delay_cnt: std_logic_vector(15 downto 0) := U16_ZERO;

signal fakesync: std_logic;
signal sync_change_cnt: std_logic_vector(15 downto 0) := U16_ZERO;


-- Buffer I/O and control signals
signal buffer_in_a: std_logic_vector(16 downto 0);
signal buffer_in_b: std_logic_vector(16 downto 0);
signal buffer_out_a: std_logic_vector(16 downto 0);
signal buffer_out_b: std_logic_vector(16 downto 0);
signal buffer_en_a: std_logic;
signal buffer_en_b: std_logic;

signal buffer_sel: std_logic; -- 0 is A, 1 is B

signal pixel_red_a: std_logic_vector(9 downto 0);
signal pixel_green_a: std_logic_vector(9 downto 0);
signal pixel_blue_a: std_logic_vector(9 downto 0);

signal pixel_red_b: std_logic_vector(9 downto 0);
signal pixel_green_b: std_logic_vector(9 downto 0);
signal pixel_blue_b: std_logic_vector(9 downto 0);

signal pixel_red_x: std_logic_vector(9 downto 0);
signal pixel_green_x: std_logic_vector(9 downto 0);
signal pixel_blue_x: std_logic_vector(9 downto 0);

signal rgb2yuv_rin: std_logic_vector(9 downto 0);
signal rgb2yuv_gin: std_logic_vector(9 downto 0);
signal rgb2yuv_bin: std_logic_vector(9 downto 0);

signal rgb2yuv_yout: std_logic_vector(9 downto 0);
signal rgb2yuv_pbout: std_logic_vector(9 downto 0);
signal rgb2yuv_prout: std_logic_vector(9 downto 0);

signal vga_hsync_buffer: std_logic;
signal vga_vsync_buffer: std_logic;

signal pixel_bus_in: std_logic_vector(16 downto 0);

signal clk_div: std_logic_vector(1 downto 0) := "00";

signal neo_pixel_concat: std_logic_vector(16 downto 0);

signal rgb2yuv_rgb_n: std_logic; -- Low for RGB mode, High for YPbPr mode
begin

	-- Both alternating line buffers
	buffer_a: entity work.linebuffer(behavioral) port map (neo_clk, buffer_en_a, buffer_in_a, buffer_out_a);
	buffer_b: entity work.linebuffer(behavioral) port map (neo_clk, buffer_en_b, buffer_in_b, buffer_out_b);

	-- Expansion from Neo-Geo pixel bus into 10-bit RGB values
	pixel_a: entity work.pixel(behavioral) port map (neo_clk, buffer_out_a, pixel_red_a, pixel_green_a, pixel_blue_a);
	pixel_b: entity work.pixel(behavioral) port map (neo_clk, buffer_out_b, pixel_red_b, pixel_green_b, pixel_blue_b);

	-- Pixel processor for pass-through 15KHz
	pixel_x: entity work.pixel(behavioral) port map (neo_clk, pixel_bus_in, pixel_red_x, pixel_green_x, pixel_blue_x);

	-- Optional YUV encoding
	rgb2yuv: entity work.rgb2yuv(behavioral) port map (rgb2yuv_rin, rgb2yuv_gin, rgb2yuv_bin, rgb2yuv_yout, rgb2yuv_pbout, rgb2yuv_prout, rgb2yuv_rgb_n);

	vga_clk <= not neo_clk;

	concatenate_pbus: process (neo_clk, neo_red, neo_green, neo_blue, neo_dak, neo_shad)
	begin
		neo_pixel_concat <= neo_red & neo_green & neo_blue & neo_dak & neo_shad;
	end process;

	clk_div_proc: process (neo_clk, fakesync_delayed)
	begin
		if (rising_edge(neo_clk)) then
			if (fakesync_delayed = '0') then
				clk_div <= "00";
			else
				clk_div <= clk_div + 1;
			end if;
		end if;
	end process;

	buffer_pixel_bus: process (neo_clk, neo_pixel_concat)
	begin
		if (rising_edge(neo_clk)) then
			if (clk_div(0) = '1') then
				if (neo_clr_n = '0') then
					pixel_bus_in <= U17_ZERO;
				else
					pixel_bus_in <= neo_pixel_concat;
				end if;
			end if;
		end if;
	end process;

	-- Output from RGB processor to DAC
	ypbpr_out: process (neo_clk, sw_ypbpr_n, rgb2yuv_prout, rgb2yuv_yout, rgb2yuv_pbout)
	begin
		-- Use the ypbpr switch to change encoding scheme
		rgb2yuv_rgb_n <= sw_ypbpr_n;
		vga_red <= rgb2yuv_prout;
		vga_green <= rgb2yuv_yout;
		vga_blue <= rgb2yuv_pbout;
	end process;

	-- Buffer selection to go to YPbPr processor
	vga_rgb_proc: process (neo_clk, sw_scanlines_n, buffer_sel, buffer_out_a, buffer_out_b)
	begin
		if (rising_edge(neo_clk)) then
			-- If we're in line doubling mode:
			if (sw_sdtv_res_n = '1') then
				-- Give the VGA inputs the processed neo-geo pixels so effects like
				-- DAK and SHAD are processed. 
				-- If 8-bit RGB is needed then just truncate the last two bits.
				if (buffer_sel = '1') then
					rgb2yuv_rin <= pixel_red_a;
					rgb2yuv_gin <= pixel_green_a;
					rgb2yuv_bin <= pixel_blue_a;
				else
					rgb2yuv_rin <= pixel_red_b;
					rgb2yuv_gin <= pixel_green_b;
					rgb2yuv_bin <= pixel_blue_b;
				end if;
			else
				-- Pass in from Neo-Geo directly
				rgb2yuv_rin <= pixel_red_x;
				rgb2yuv_gin <= pixel_green_x;
				rgb2yuv_bin <= pixel_blue_x;
			end if;
		end if;	
	end process;

	-- Set VGA sync stuff
	vga_sync_out: process (neo_clk)
	begin
		if (rising_edge(neo_clk)) then
			vga_hsync <= vga_hsync_buffer;
			vga_vsync <= vga_vsync_buffer;
		end if;
	end process;

	-- VGA output horizontal sync and blanking
	vga_hsync_proc: process (neo_clk, vga_pxcount, line_count, sw_ypbpr_n)
	begin
		if (rising_edge(neo_clk)) then
			-- If we're in line doubling mode:
			if (sw_sdtv_res_n = '1') then
				-- Two hsyncs for every 1 neo-geo hsync
				if (vga_pxcount >= VGA_HSYNC_START and vga_pxcount < VGA_HSYNC_END) then
					vga_hsync_buffer <= '0';
				else
					vga_hsync_buffer <= '1';
				end if;
				
				-- Shouldn't really be needed since the image in the line buffers 
				-- has blanking of its own, but it is safer to blank it here too.
				if ((vga_pxcount >= VGA_VISIBLE_START and vga_pxcount < VGA_VISIBLE_END) or sw_ypbpr_n = '0') then
					vga_blank <= '1';
				else
					vga_blank <= '0';
				end if;
			-- For 15Khz output
			else
				-- Pass timings unchanged. Hsync pin is used for C-sync with the VGA connector.
				vga_hsync_buffer <= neo_csync;
				
				if (sw_ypbpr_n = '1') then
					vga_blank <= neo_clr_n;
				else
					-- In YpbPr, we avoid the blanking pin as it malforms the sync signal.
					vga_blank <= '1';
				end if;
			end if;
		end if;
	end process;

	vga_csync_out: process (neo_clk, sw_ypbpr_n)
	begin
		if (rising_edge(neo_clk)) then
			if (sw_ypbpr_n = '0' or j_want_sog_n = '0') then -- Sync on green/Y is only for YpbPr, or when forced
				if (sw_sdtv_res_n = '1') then
					-- Generate composite sync for the Y channel / Sync-on-green
					vga_sync <= vga_hsync_buffer xnor vga_vsync_buffer;
				else
					-- Pass through the Neo-Geo's composite sync to exactly match original timings
					vga_sync <= neo_csync;
				end if;
			else
				-- In RGB mode, no sync is injected into the green output
				vga_sync <= '0';
			end if;
		end if;
	end process;

	-- VGA output vertical sync
	vga_vsync_proc: process (neo_clk, vsync_count, line_count)
	begin
		if (rising_edge(neo_clk)) then
			if (line_count >= VGA_VSYNC_LINE_START and line_count < VGA_VSYNC_LINE_END) then
				vga_vsync_buffer <= '0';
			else
				vga_vsync_buffer <= '1';
			end if;
		end if;
	end process;


	-- Control pixel count and buffer alternation
	pixel_inc: process(neo_clk, neo_pxcount, vsync_count)
	begin
		if (rising_edge(neo_clk)) then
			if (sw_sdtv_res_n = '1') then
				-- Process vsync two lines after the Neo does it so the buffer swap
				-- doesn't stop until after the last line.
				-- This is what keeps the image synchronized (and thus centered)
				if (vsync_count = (NEO_LINE_LEN * 2)) then
					line_count <= U16_ZERO;
					neo_pxcount <= U16_ZERO;
				elsif (neo_pxcount = (NEO_LINE_LEN - 1)) then
					-- End of Neo-Geo line. Swap buffers
					buffer_sel <= not buffer_sel;
					-- Bottom of screen, reset line count
					if (line_count = NUM_LINES) then
						line_count <= U16_ZERO;
					else
						line_count <= line_count + 1;
					end if;
					neo_pxcount <= U16_ZERO;
				else
					neo_pxcount <= neo_pxcount + 1;
				end if;
				
				if (vsync_count = NEO_LINE_LEN) then
					vga_pxcount <= U16_ZERO;
				elsif (vga_pxcount = VGA_LINE_LEN - 1) then
					vga_pxcount <= U16_ZERO;
				else
					vga_pxcount <= vga_pxcount + 1;
				end if;
			end if;
		end if;
	end process;

	-- Detect if the system is a NEO-GRZ based system, and change H-Shift as needed
	detect_grz: process(neo_clk, neo_clr_n)
	begin
		if (rising_edge(neo_clk)) then	
			--if (line_count = 16 and neo_clr_n = '0') then -- Only the NEO-GRZ blanks horizontally.
			--	h_shift <= NEO_GRZ_SHIFT;
			--end if;
			if (j_mv1c_sel_n = '0') then
				h_shift <= NEO_GRZ_SHIFT;
			else
				h_shift <= NEO_B1_SHIFT;
			end if;
		end if;
	end process;	

	-- Generate a fake VSync signal from the Neo-Geo's CSync
	make_fakesync: process(neo_clk, neo_csync)
	begin
		if (rising_edge(neo_clk)) then
			if (neo_csync /= fakesync) then
				-- The change must be observed for greater than the threshhold before it "sticks".
				-- This is a crude 1-bit-resolution low pass filter with an exact cutoff. 
				if (sync_change_cnt >= FAKESYNC_THRESH) then
					fakesync <= neo_csync;
				else
					sync_change_cnt <= sync_change_cnt + 1;
				end if;
			else
				sync_change_cnt <= U16_ZERO;
			end if;
			
			-- Show the interpreted VSync signal as an indicator that the system is operating correctly. 
			led_out <= not fakesync;		
		end if;
	end process;

	-- Make a delayed sync
	make_delayed_sync: process(neo_clk, fakesync)
	begin
		if (rising_edge(neo_clk)) then
			if (fakesync /= fakesync_delayed) then
				if (sync_delay_cnt >= h_shift) then
					fakesync_delayed <= neo_csync;
				else
					sync_delay_cnt <= sync_delay_cnt + 1;
				end if;
			else
				sync_delay_cnt <= U16_ZERO;
			end if;
		end if;
	end process;

	-- Count how long Vsync has been active on the Neo-Geo
	vsync_counter: process(neo_clk, fakesync_delayed)
	begin
		if (rising_edge(neo_clk)) then
			if (fakesync_delayed = '0') then
				vsync_count <= vsync_count + 1;
			else
				vsync_count <= U16_ZERO;
			end if;
		end if;
	end process;

	-- Manage capturing and buffer input prouting
	capture_data: process(neo_clk, buffer_sel, sw_scanlines_n)
	begin
		if (rising_edge(neo_clk)) then
			if (sw_sdtv_res_n = '1') then
				if (buffer_sel = '0') then
					-- Concatenate Neo-Geo pixel bus into a single "pixel" vector
					if (line_count < NUM_LINES-1 and neo_clr_n = '1') then
						buffer_in_a <= neo_pixel_concat;
					else
						buffer_in_a <= U17_ZERO;
					end if;
				
					-- Capture on every other double-pixel-clock
					buffer_en_a <= neo_pxcount(0);
					
					if (sw_scanlines_n(1) = '0') then -- Full dark scanlines
						buffer_in_b <= U17_ZERO;
					elsif (sw_scanlines_n(0) = '0') then -- Partially darkened scanlines
						buffer_in_b <= '0' & buffer_out_b(16 downto 13) & '0' & buffer_out_b(11 downto 8) & '0' & buffer_out_b(6 downto 3) & "00";
					else
						buffer_in_b <= buffer_out_b; -- No scanlines
					end if;
					
					-- Shift out other buffer full- speed for VGA output
					buffer_en_b <= '1';
				else
					-- Concatenate Neo-Geo pixel bus into a single 'pixel' vector
					if (line_count < NUM_LINES-1 and neo_clr_n = '1') then
						buffer_in_b <= neo_pixel_concat;
					else
						buffer_in_b <= U17_ZERO;
					end if;

					-- Capture on every other double-pixel-clock
					buffer_en_b <= neo_pxcount(0);
					
					if (sw_scanlines_n(1) = '0') then
						buffer_in_a <= U17_ZERO;
					elsif (sw_scanlines_n(0) = '0') then
						buffer_in_a <= '0' & buffer_out_a(16 downto 13) & '0' & buffer_out_a(11 downto 8) & '0' & buffer_out_a(6 downto 3) & "00";
					else
						buffer_in_a <= buffer_out_a;
					end if;

					-- Shift out other buffer full- speed for VGA output
					buffer_en_a <= '1';
				end if;
			end if;
		end if;
	end process;
end behavioral;
